/*
    https://hdlbits.01xz.net/wiki/Module_cseladd
*/

module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    wire [15:0] sum1, sum2, sum3, sum_sel;
    wire cout1, cout2, cout3;

    add16 inst1 (.a(a[15:0]), .b(b[15:0]), .cin(0), .sum(sum1), .cout(cout1));
    add16 inst2 (.a(a[31:16]), .b(b[31:16]), .cin(0), .sum(sum2), .cout(cout2));
    add16 inst3 (.a(a[31:16]), .b(b[31:16]), .cin(1), .sum(sum3), .cout(cout3));

    assign sum_sel = cout1 ? sum3 : sum2;
    assign sum = {sum_sel, sum1};

endmodule

module add16 ( input[15:0] a, input[15:0] b, input cin, output[15:0] sum, output cout );
endmodule
